// Description
// ### Author : Md Nazmus Sakib(email)

`include "config_pkg.sv"
//`include "axi4l_assign.svh"
//`include "axi4l_typedef.svh"
//`include "axi4_assign.svh"
//`include "axi4_typedef.svh"
//`include "default_param_pkg.sv"

import config_pkg::uinstr_t;
import config_pkg::data_t;
import config_pkg::w_data_t;
import config_pkg::code_t;
module receive_fsm(
    input logic clk,
    input logic arst_ni,
    input logic rd_data_valid_i,
    input data_t rd_data_i,
    output data_t operand_a_o,
    output data_t operand_b_o,
    output w_data_t operand_c_o,
    output logic operation_valid_o
  );

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////

  typedef enum logic [1:0] {oper_a, oper_b, oper_c, oper_c_2} State;
  State currentstate, nextstate;
  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////
  data_t reg_a;
  data_t reg_b;
  data_t reg_c;
  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////




  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIAL{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////
  always_ff @(posedge clk)
  begin
    if (~arst_ni)
    begin
      currentstate <= oper_a;
    end
    else
    begin
      currentstate <= nextstate;
    end
  end
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-Combinational{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //State Assignment


  always_comb
  begin
    operand_a_o = 0;
    operand_b_o = 0;
    operand_c_o = 0;
    operation_valid_o =0;
    case (currentstate)
      oper_a:
      begin
        if (rd_data_valid_i)
        begin
          reg_a = rd_data_i;
          operation_valid_o =0;
          nextstate = oper_b;
        end
        else
          nextstate = oper_a;
      end

      oper_b:
      begin
        if (rd_data_valid_i)
        begin
          reg_b = rd_data_i;
          nextstate = oper_c;
        end
        else
          nextstate = oper_b;
      end

      oper_c:
      begin
        if (rd_data_valid_i)
        begin
          reg_c = rd_data_i;
          nextstate = oper_c_2;
        end
        else
          nextstate = oper_c;
      end

      oper_c_2:
      begin
        if (rd_data_valid_i)
        begin
          operand_a_o = reg_a;
          operand_b_o = reg_b;
          operand_c_o = {reg_c, rd_data_i};
          operation_valid_o =1;
          nextstate = oper_a;
        end
        else
          nextstate = oper_c_2;
      end
    endcase
  end
endmodule
