`define ADDR_MATCHING(__HSUINSTR__, __SRC_CLK__, __DEST_CLK__) 
  bit Fail = 0;
